
// apb_pkg

package apb_pkg;

// include/import necessary files here





endpackage : apb_pkg
